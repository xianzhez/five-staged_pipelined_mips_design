library verilog;
use verilog.vl_types.all;
entity top_tb_v is
end top_tb_v;
