library verilog;
use verilog.vl_types.all;
entity Decode is
    generic(
        R_type_op       : integer := 0;
        ADD_funct       : integer := 32;
        ADDU_funct      : integer := 33;
        AND_funct       : integer := 36;
        XOR_funct       : integer := 38;
        OR_funct        : integer := 37;
        NOR_funct       : integer := 39;
        SUB_funct       : integer := 34;
        SUBU_funct      : integer := 35;
        SLT_funct       : integer := 42;
        SLTU_funct      : integer := 43;
        SLL_funct       : integer := 0;
        SLLV_funct      : integer := 4;
        SRL_funct       : integer := 2;
        SRLV_funct      : integer := 6;
        SRA_funct       : integer := 3;
        SRAV_funct      : integer := 7;
        JR_funct        : integer := 8;
        BEQ_op          : integer := 4;
        BNE_op          : integer := 5;
        BGEZ_op         : integer := 1;
        BGEZ_rt         : integer := 1;
        BGTZ_op         : integer := 7;
        BGTZ_rt         : integer := 0;
        BLEZ_op         : integer := 6;
        BLEZ_rt         : integer := 0;
        BLTZ_op         : integer := 1;
        BLTZ_rt         : integer := 0;
        J_op            : integer := 2;
        ADDI_op         : integer := 8;
        ADDIU_op        : integer := 9;
        ANDI_op         : integer := 12;
        XORI_op         : integer := 14;
        ORI_op          : integer := 13;
        SLTI_op         : integer := 10;
        SLTIU_op        : integer := 11;
        SW_op           : integer := 43;
        LW_op           : integer := 35;
        alu_add         : integer := 0;
        alu_and         : integer := 1;
        alu_xor         : integer := 2;
        alu_or          : integer := 3;
        alu_nor         : integer := 4;
        alu_sub         : integer := 5;
        alu_andi        : integer := 6;
        alu_xori        : integer := 7;
        alu_ori         : integer := 8;
        alu_jr          : integer := 9;
        alu_beq         : integer := 10;
        alu_bne         : integer := 11;
        alu_bgez        : integer := 12;
        alu_bgtz        : integer := 13;
        alu_blez        : integer := 14;
        alu_bltz        : integer := 15;
        alu_sll         : integer := 16;
        alu_srl         : integer := 17;
        alu_sra         : integer := 18;
        alu_slt         : integer := 19;
        alu_sltu        : integer := 20
    );
    port(
        MemtoReg        : out    vl_logic;
        RegWrite        : out    vl_logic;
        MemWrite        : out    vl_logic;
        MemRead         : out    vl_logic;
        ALUCode         : out    vl_logic_vector(4 downto 0);
        ALUSrcA         : out    vl_logic;
        ALUSrcB         : out    vl_logic;
        RegDst          : out    vl_logic;
        J               : out    vl_logic;
        JR              : out    vl_logic;
        Instruction     : in     vl_logic_vector(31 downto 0)
    );
end Decode;
